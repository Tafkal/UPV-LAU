LIBRARY ieee;
USE ieee.std_logic_1164.all;

package Q_val is
	constant Q : integer := 10;
end Q_val;